library verilog;
use verilog.vl_types.all;
entity test_block_vlg_vec_tst is
end test_block_vlg_vec_tst;
